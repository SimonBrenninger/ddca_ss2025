
entity util_tb is
end entity;

architecture test of util_tb is 
begin

end architecture;



