library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.vga_ctrl_pkg.all;


architecture arch of vga_ctrl is
	-- TODO: Add signals, constants, types and subprograms as needed
begin

	-- TODO: Implement the vga_ctrl

end architecture;


