library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.snes_ctrl_pkg.all;


architecture arch of snes_ctrl is
	-- TODO: Declare signals, subprograms, constants and types as needed
begin

	-- TODO: Implement

end architecture;
