library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.sorting_network_pkg.all;

architecture arch_combinatorial of sorting_network is

begin

end architecture;
