
library ieee;
use ieee.std_logic_1164.all;
use work.gfx_core_pkg.all;

package gfx_init_pkg is
	type gfx_init_cmds_t is array(natural range<>) of gfx_cmd_t;

	constant GFX_INIT_CMDS : gfx_init_cmds_t(0 to 2783) := (
		x"9000",
		x"0000",
		x"0000",
		x"0140",
		x"00f0",
		x"9001",
		x"2c00",
		x"0001",
		x"0140",
		x"00f0",
		x"9002",
		x"5800",
		x"0002",
		x"0158",
		x"0008",
		x"7001",
		x"0560",
		x"5800",
		x"0002",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"0000",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"00ff",
		x"ff00",
		x"ffff",
		x"0000",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"0000",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"ff00",
		x"0000",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"0000",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"9003",
		x"62c0",
		x"0002",
		x"00c0",
		x"000c",
		x"7001",
		x"0480",
		x"62c0",
		x"0002",
		x"2424",
		x"2424",
		x"2424",
		x"2424",
		x"2424",
		x"2424",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"4900",
		x"0049",
		x"0000",
		x"0000",
		x"4900",
		x"0049",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"006d",
		x"6d6d",
		x"6d6d",
		x"006d",
		x"9292",
		x"0000",
		x"0000",
		x"0000",
		x"2424",
		x"2524",
		x"2525",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"4924",
		x"926d",
		x"6d92",
		x"6d6d",
		x"6d6d",
		x"246d",
		x"b66d",
		x"92b6",
		x"9292",
		x"9292",
		x"b692",
		x"6db6",
		x"4949",
		x"6d00",
		x"006d",
		x"6d00",
		x"006d",
		x"4949",
		x"db00",
		x"dbdb",
		x"dbdb",
		x"dbdb",
		x"dbdb",
		x"00db",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"db00",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"00db",
		x"6d6d",
		x"db6d",
		x"6d6d",
		x"6d6d",
		x"6ddb",
		x"6d6d",
		x"ff6d",
		x"dbdb",
		x"00db",
		x"db00",
		x"dbdb",
		x"6dff",
		x"6d6d",
		x"006d",
		x"6d92",
		x"6d6d",
		x"006d",
		x"6d92",
		x"0000",
		x"0000",
		x"0000",
		x"2424",
		x"2524",
		x"2525",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"00ff",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"6d24",
		x"b692",
		x"b6b6",
		x"b6b6",
		x"92b6",
		x"246d",
		x"b66d",
		x"4992",
		x"926d",
		x"6d92",
		x"9249",
		x"6db6",
		x"0049",
		x"6d6d",
		x"b600",
		x"00b6",
		x"6d6d",
		x"4900",
		x"db00",
		x"b6b6",
		x"b6b6",
		x"b6b6",
		x"b6b6",
		x"00db",
		x"4949",
		x"6d6d",
		x"496d",
		x"6d49",
		x"6d6d",
		x"4949",
		x"6d00",
		x"dbdb",
		x"4949",
		x"4949",
		x"dbdb",
		x"006d",
		x"db6d",
		x"db6d",
		x"006d",
		x"6d00",
		x"6ddb",
		x"6ddb",
		x"db6d",
		x"ffda",
		x"2449",
		x"4924",
		x"daff",
		x"6ddb",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"2424",
		x"2524",
		x"2525",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"00ff",
		x"6d24",
		x"b692",
		x"b6b6",
		x"b6b6",
		x"92b6",
		x"246d",
		x"926d",
		x"246d",
		x"9225",
		x"2592",
		x"6d24",
		x"6d92",
		x"6d00",
		x"006d",
		x"b6b6",
		x"b6b6",
		x"6d00",
		x"006d",
		x"db00",
		x"00b6",
		x"0000",
		x"0000",
		x"b600",
		x"00db",
		x"4949",
		x"6d6d",
		x"496d",
		x"6d49",
		x"6d6d",
		x"4949",
		x"6d00",
		x"dbdb",
		x"4949",
		x"4949",
		x"dbdb",
		x"006d",
		x"db6d",
		x"6d6d",
		x"006d",
		x"6d00",
		x"6d6d",
		x"6ddb",
		x"b66d",
		x"24ff",
		x"6d24",
		x"246d",
		x"ff24",
		x"6db6",
		x"9292",
		x"6d6d",
		x"006d",
		x"9292",
		x"6d6d",
		x"006d",
		x"4949",
		x"4949",
		x"4949",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"0000",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"00ff",
		x"6d24",
		x"b6b6",
		x"b6b6",
		x"dbb6",
		x"b6b6",
		x"2492",
		x"b66d",
		x"4992",
		x"926d",
		x"6d92",
		x"9249",
		x"6db6",
		x"6d00",
		x"b600",
		x"00b6",
		x"b600",
		x"00b6",
		x"006d",
		x"db00",
		x"00b6",
		x"4949",
		x"4949",
		x"b600",
		x"00db",
		x"6d49",
		x"6d49",
		x"db49",
		x"49db",
		x"496d",
		x"496d",
		x"6d00",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"006d",
		x"db6d",
		x"6ddb",
		x"0000",
		x"0000",
		x"db6d",
		x"6ddb",
		x"ff6d",
		x"0049",
		x"6d49",
		x"496d",
		x"4900",
		x"6dff",
		x"6d92",
		x"6d6d",
		x"006d",
		x"6d92",
		x"6d6d",
		x"006d",
		x"4949",
		x"4949",
		x"4949",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"00ff",
		x"6d24",
		x"b692",
		x"dbb6",
		x"dbdb",
		x"b6b6",
		x"2492",
		x"b66d",
		x"b6b6",
		x"92b6",
		x"b692",
		x"b6b6",
		x"6db6",
		x"0000",
		x"b6b6",
		x"b600",
		x"00b6",
		x"b6b6",
		x"0000",
		x"db00",
		x"00b6",
		x"4949",
		x"4949",
		x"b600",
		x"00db",
		x"4949",
		x"496d",
		x"dbdb",
		x"dbdb",
		x"6d49",
		x"4949",
		x"6d00",
		x"4949",
		x"db49",
		x"49db",
		x"4949",
		x"006d",
		x"006d",
		x"6ddb",
		x"6d00",
		x"006d",
		x"db6d",
		x"6d00",
		x"006d",
		x"6d00",
		x"6d6d",
		x"6d6d",
		x"006d",
		x"6d00",
		x"6d92",
		x"6d6d",
		x"006d",
		x"6d92",
		x"6d6d",
		x"006d",
		x"4949",
		x"4949",
		x"4949",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"6d24",
		x"b692",
		x"dbb6",
		x"dbdb",
		x"92b6",
		x"246d",
		x"b66d",
		x"b6b6",
		x"92b6",
		x"b692",
		x"b6b6",
		x"6db6",
		x"0000",
		x"b6b6",
		x"b600",
		x"00b6",
		x"b6b6",
		x"0000",
		x"db00",
		x"00b6",
		x"4949",
		x"4949",
		x"b600",
		x"00db",
		x"4949",
		x"496d",
		x"dbdb",
		x"dbdb",
		x"6d49",
		x"4949",
		x"6d00",
		x"4949",
		x"db49",
		x"49db",
		x"4949",
		x"006d",
		x"6d00",
		x"00db",
		x"006d",
		x"6d00",
		x"db00",
		x"006d",
		x"006d",
		x"6d00",
		x"6d6d",
		x"6d6d",
		x"006d",
		x"6d00",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"9292",
		x"9292",
		x"9292",
		x"b6b6",
		x"b6b6",
		x"b6b6",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"00ff",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"6d24",
		x"b692",
		x"b6b6",
		x"b6db",
		x"92b6",
		x"246d",
		x"b66d",
		x"4992",
		x"926d",
		x"6d92",
		x"9249",
		x"6db6",
		x"6d00",
		x"b600",
		x"00b6",
		x"b600",
		x"00b6",
		x"006d",
		x"db00",
		x"00b6",
		x"4949",
		x"4949",
		x"b600",
		x"00db",
		x"6d49",
		x"6d49",
		x"db49",
		x"49db",
		x"496d",
		x"496d",
		x"6d00",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"006d",
		x"db00",
		x"00db",
		x"6d6d",
		x"6d6d",
		x"db00",
		x"00db",
		x"ff6d",
		x"0049",
		x"6d49",
		x"496d",
		x"4900",
		x"6dff",
		x"006d",
		x"9292",
		x"6d6d",
		x"006d",
		x"9292",
		x"6d6d",
		x"9292",
		x"9292",
		x"9292",
		x"b6b6",
		x"b6b6",
		x"b6b6",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"ffff",
		x"00ff",
		x"0000",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"00ff",
		x"6d24",
		x"b692",
		x"b6b6",
		x"b6b6",
		x"b6b6",
		x"2492",
		x"926d",
		x"246d",
		x"9225",
		x"2592",
		x"6d24",
		x"6d92",
		x"6d00",
		x"006d",
		x"b6b6",
		x"b6b6",
		x"6d00",
		x"006d",
		x"db00",
		x"00b6",
		x"0000",
		x"0000",
		x"b600",
		x"00db",
		x"4949",
		x"6d6d",
		x"496d",
		x"6d49",
		x"6d6d",
		x"4949",
		x"6d00",
		x"dbdb",
		x"4949",
		x"4949",
		x"dbdb",
		x"006d",
		x"db00",
		x"0000",
		x"6d00",
		x"006d",
		x"0000",
		x"00db",
		x"b66d",
		x"24ff",
		x"6d24",
		x"246d",
		x"ff24",
		x"6db6",
		x"006d",
		x"6d92",
		x"6d6d",
		x"006d",
		x"6d92",
		x"6d6d",
		x"9292",
		x"9292",
		x"9292",
		x"b6b6",
		x"b6b6",
		x"b6b6",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"00ff",
		x"6d24",
		x"b6b6",
		x"b6b6",
		x"b6b6",
		x"92b6",
		x"246d",
		x"b66d",
		x"4992",
		x"926d",
		x"6d92",
		x"9249",
		x"6db6",
		x"0049",
		x"6d6d",
		x"b600",
		x"00b6",
		x"6d6d",
		x"4900",
		x"db00",
		x"b6b6",
		x"b6b6",
		x"b6b6",
		x"b6b6",
		x"00db",
		x"4949",
		x"6d6d",
		x"496d",
		x"6d49",
		x"6d6d",
		x"4949",
		x"6d00",
		x"dbdb",
		x"4949",
		x"4949",
		x"dbdb",
		x"006d",
		x"db00",
		x"db00",
		x"6d00",
		x"006d",
		x"00db",
		x"00db",
		x"db6d",
		x"ffda",
		x"2449",
		x"4924",
		x"daff",
		x"6ddb",
		x"006d",
		x"6d92",
		x"6d6d",
		x"006d",
		x"6d92",
		x"6d6d",
		x"dada",
		x"dbda",
		x"dbdb",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"00ff",
		x"6d24",
		x"b692",
		x"92b6",
		x"92b6",
		x"9292",
		x"246d",
		x"b66d",
		x"92b6",
		x"9292",
		x"9292",
		x"b692",
		x"6db6",
		x"4949",
		x"6d00",
		x"006d",
		x"6d00",
		x"006d",
		x"4949",
		x"db00",
		x"dbdb",
		x"dbdb",
		x"dbdb",
		x"dbdb",
		x"00db",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"db00",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"00db",
		x"0000",
		x"db00",
		x"0000",
		x"0000",
		x"00db",
		x"0000",
		x"ff6d",
		x"dbdb",
		x"00db",
		x"db00",
		x"dbdb",
		x"6dff",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"dada",
		x"dbda",
		x"dbdb",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ff00",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ff00",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"ff00",
		x"ffff",
		x"00ff",
		x"0000",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"2424",
		x"2424",
		x"2424",
		x"2424",
		x"2424",
		x"2424",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"4900",
		x"0049",
		x"0000",
		x"0000",
		x"4900",
		x"0049",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"4949",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d6d",
		x"6d92",
		x"006d",
		x"9292",
		x"6d6d",
		x"006d",
		x"9292",
		x"dada",
		x"dbda",
		x"dbdb",
		x"ffff",
		x"ffff",
		x"ffff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"00ff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"ffff",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"0000",
		x"807a",
		x"80d8",
		x"80c5",
		x"802c",
		x"809e",
		x"80bc",
		x"8006",
		x"8044",
		x"80d0",
		x"80fc",
		x"8010",
		x"8058",
		x"80d6",
		x"80cd",
		x"803b",
		x"80c6",
		x"805f",
		x"80df",
		x"8018",
		x"80ea",
		x"8085",
		x"80ae",
		x"8030",
		x"808b",
		x"8085",
		x"801e",
		x"807b",
		x"8003",
		x"8066",
		x"8034",
		x"80b5",
		x"808b",
		x"80cf",
		x"800c",
		x"80dd",
		x"80f2",
		x"80e5",
		x"80e6",
		x"808c",
		x"8001",
		x"8002",
		x"80cb",
		x"8022",
		x"80d4",
		x"809b",
		x"802c",
		x"80df",
		x"80b7",
		x"809e",
		x"80e3",
		x"80ad",
		x"8080",
		x"8012",
		x"805e",
		x"8061",
		x"8089",
		x"8085",
		x"8033",
		x"8045",
		x"80d7",
		x"8057",
		x"80fd",
		x"8030",
		x"8016",
		x"8068",
		x"80f3",
		x"80bb",
		x"8035",
		x"80dc",
		x"80fe",
		x"8076",
		x"8017",
		x"80a5",
		x"8020",
		x"8007",
		x"803a",
		x"80ba",
		x"80a1",
		x"80b0",
		x"8091",
		x"80dd",
		x"8078",
		x"807c",
		x"80ca",
		x"800e",
		x"8034",
		x"800f",
		x"801b",
		x"802e",
		x"8060",
		x"8065",
		x"80ce",
		x"80df",
		x"80b6",
		x"8001",
		x"80c2",
		x"8033",
		x"8002",
		x"8010",
		x"80b3",
		x"808a",
		x"802d",
		x"800e",
		x"80b1",
		x"8065",
		x"80bd",
		x"80be",
		x"8003",
		x"80b6",
		x"8023",
		x"80e5",
		x"80c1",
		x"8056",
		x"8034",
		x"8069",
		x"80e7",
		x"8067",
		x"80b9",
		x"8051",
		x"8089",
		x"8079",
		x"8091",
		x"80e8",
		x"8031",
		x"802e",
		x"806a",
		x"80c9",
		x"8029",
		x"8065",
		x"8059",
		x"8065",
		x"80d0",
		x"80a5",
		x"8073",
		x"8062",
		x"8060",
		x"80fd",
		x"8004",
		x"8027",
		x"80d1",
		x"8080",
		x"80c4",
		x"806b",
		x"8069",
		x"9007",
		x"6bc0",
		x"0002",
		x"000c",
		x"000c",
		x"7001",
		x"0048",
		x"6bc0",
		x"0002",
		x"f152",
		x"04e5",
		x"9cb7",
		x"6d2e",
		x"d4f0",
		x"7839",
		x"a582",
		x"e65e",
		x"b639",
		x"996a",
		x"8ef1",
		x"ee40",
		x"6df7",
		x"6d14",
		x"4346",
		x"e4dd",
		x"7fef",
		x"9cb8",
		x"9581",
		x"60ac",
		x"a322",
		x"ba43",
		x"01ff",
		x"c5bb",
		x"94ff",
		x"a0c3",
		x"3762",
		x"fd02",
		x"41f0",
		x"f720",
		x"9b38",
		x"7710",
		x"d306",
		x"54de",
		x"8aaf",
		x"6513",
		x"4585",
		x"5d60",
		x"d59a",
		x"b1df",
		x"1cb9",
		x"ab1f",
		x"514e",
		x"686c",
		x"1400",
		x"b910",
		x"d3b6",
		x"ec6f",
		x"6152",
		x"d23e",
		x"0dfe",
		x"d879",
		x"d109",
		x"619e",
		x"03d3",
		x"b684",
		x"4637",
		x"820d",
		x"9903",
		x"a930",
		x"fe1b",
		x"4486",
		x"4a5d",
		x"46b9",
		x"370c",
		x"fe11",
		x"5b85",
		x"404b",
		x"2dd5",
		x"f907",
		x"e4a9",
		x"4043",
		x"9800",
		x"80ff",
		x"8400"
	);
end package;

