library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.gc_ctrl_pkg.all;

architecture arch of gc_ctrl is

	-- TODO: Declare signals, subprograms, constants and types as needed

begin

	-- TODO: Implement

end architecture;
